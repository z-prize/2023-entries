`define SHADD_6(_W, _O, _S0, _S1, _S2, _S3, _S4, _S5, _I0, _I1, _I2, _I3, _I4, _I5) shift_adder_6 #(.W(_W),.S0(_S0),.S1(_S1),.S2(_S2),.S3(_S3),.S4(_S4),.S5(_S5),.R(1)) ``_O``_shadd6_inst (.in0(_I0),.in1(_I1),.in2(_I2),.in3(_I3),.in4(_I4),.in5(_I5),.out0(_O),.clk(clk),.rst(rst));

module zprize_mul_384_shift #(
    W=384,W0=W,W1=W,L=3,T=32'h07F7_F999,
    W2=W/2,
    R_I=0,
    CT = T[0 +: 4],
    ST = T >> 4,
    M=32,
    S=0
)(
    input wire                                                      clk,
    input wire                                                      rst,

    input wire [W0-1:0]                                             in0,
    input wire [W1-1:0]                                             in1,
    input wire [M-1:0]                                              m_i,
    output logic [M-1:0]                                            m_o,
    output logic [W0+W1-1:0]                                        out0
);

logic [W0-1:0] in0_r;
logic [W1-1:0] in1_r;
logic [M-1:0] m_i_r;

//////////////////////////////////////////////////////////////////////////////
///////////////////////    RTL BODY        ///////////////////////////////////
//////////////////////////////////////////////////////////////////////////////

        assign in0_r = in0;
        assign in1_r = in1;
        assign m_i_r = m_i;


logic [384-1:0] out_p;
logic [384-1:0] out_n;
logic [M-1:0] p_m_o;
logic [M-1:0] n_m_o;
logic [6-1:0][M-1:0] p_m_o_p;
logic [164-1:0] p_s_0_24;
logic [ 90-1:0] p_s_0_36;
logic [ 90-1:0] p_s_1_06;
logic [336-1:0] p_s_1_00;
logic [ 11-1:0] p_s_0_48;
logic [120-1:0] p_s_0_30;
logic [ 50-1:0] p_s_0_42;
logic [208-1:0] p_s_0_18;
logic [336-1:0] p_s_2_00;
logic [336-1:0] p_s_0_00;
logic [277-1:0] p_s_0_06;
logic [236-1:0] p_s_0_12;
`SHADD_6(336, p_s_0_00,   0,   3,   8,  10,  15,  45, {336'b0, in0[0+:336]}, {336'b0, in0[0+:333]}, {336'b0, in0[0+:328]}, {336'b0, in0[0+:326]}, {336'b0, in0[0+:321]}, {336'b0, in0[0+:291]});
`SHADD_6(277, p_s_0_06,   0,   3,   5,   8,  14,  17, {277'b0, in0[0+:277]}, {277'b0, in0[0+:274]}, {277'b0, in0[0+:272]}, {277'b0, in0[0+:269]}, {277'b0, in0[0+:263]}, {277'b0, in0[0+:260]});
`SHADD_6(236, p_s_0_12,   0,   9,  15,  18,  22,  24, {236'b0, in0[0+:236]}, {236'b0, in0[0+:227]}, {236'b0, in0[0+:221]}, {236'b0, in0[0+:218]}, {236'b0, in0[0+:214]}, {236'b0, in0[0+:212]});
`SHADD_6(208, p_s_0_18,   0,  14,  18,  20,  25,  40, {208'b0, in0[0+:208]}, {208'b0, in0[0+:194]}, {208'b0, in0[0+:190]}, {208'b0, in0[0+:188]}, {208'b0, in0[0+:183]}, {208'b0, in0[0+:168]});
`SHADD_6(164, p_s_0_24,   0,   7,  19,  22,  25,  35, {164'b0, in0[0+:164]}, {164'b0, in0[0+:157]}, {164'b0, in0[0+:145]}, {164'b0, in0[0+:142]}, {164'b0, in0[0+:139]}, {164'b0, in0[0+:129]});
`SHADD_6(120, p_s_0_30,   0,   6,   9,  11,  15,  25, {120'b0, in0[0+:120]}, {120'b0, in0[0+:114]}, {120'b0, in0[0+:111]}, {120'b0, in0[0+:109]}, {120'b0, in0[0+:105]}, {120'b0, in0[0+: 95]});
`SHADD_6( 90, p_s_0_36,   0,   2,  20,  23,  26,  32, {90'b0, in0[0+: 90]}, {90'b0, in0[0+: 88]}, {90'b0, in0[0+: 70]}, {90'b0, in0[0+: 67]}, {90'b0, in0[0+: 64]}, {90'b0, in0[0+: 58]});
`SHADD_6( 50, p_s_0_42,   0,   5,  25,  31,  34,  36, {50'b0, in0[0+: 50]}, {50'b0, in0[0+: 45]}, {50'b0, in0[0+: 25]}, {50'b0, in0[0+: 19]}, {50'b0, in0[0+: 16]}, {50'b0, in0[0+: 14]});
`SHADD_6( 11, p_s_0_48,   0,   0,   0,   0,   0,   0, {11'b0, in0[0+: 11]}, {11'b0, '0}, {11'b0, '0}, {11'b0, '0}, {11'b0, '0}, {11'b0, '0});
`SHADD_6(336, p_s_1_00,   0,  59, 100, 128, 172, 216, {336'b0, p_s_0_00}, {336'b0, p_s_0_06}, {336'b0, p_s_0_12}, {336'b0, p_s_0_18}, {336'b0, p_s_0_24}, {336'b0, p_s_0_30});
`SHADD_6( 90, p_s_1_06,   0,  40,  79,   0,   0,   0, {90'b0, p_s_0_36}, {90'b0, p_s_0_42}, {90'b0, p_s_0_48}, {90'b0, '0}, {90'b0, '0}, {90'b0, '0});
`SHADD_6(336, p_s_2_00,   0, 246,   0,   0,   0,   0, {336'b0, p_s_1_00}, {336'b0, p_s_1_06}, {336'b0, '0}, {336'b0, '0}, {336'b0, '0}, {336'b0, '0});
assign out_p = p_s_2_00 << 48;
assign p_m_o = p_m_o_p[6-1];
always@(posedge clk) p_m_o_p[0] <= m_i;
always@(posedge clk) p_m_o_p[1] <= p_m_o_p[1-1];
always@(posedge clk) p_m_o_p[2] <= p_m_o_p[2-1];
always@(posedge clk) p_m_o_p[3] <= p_m_o_p[3-1];
always@(posedge clk) p_m_o_p[4] <= p_m_o_p[4-1];
always@(posedge clk) p_m_o_p[5] <= p_m_o_p[5-1];
logic [6-1:0][M-1:0] n_m_o_p;
logic [107-1:0] n_s_0_36;
logic [136-1:0] n_s_0_30;
logic [166-1:0] n_s_0_24;
logic [  2-1:0] n_s_0_48;
logic [267-1:0] n_s_0_06;
logic [384-1:0] n_s_0_00;
logic [229-1:0] n_s_0_12;
logic [107-1:0] n_s_1_06;
logic [ 52-1:0] n_s_0_42;
logic [384-1:0] n_s_1_00;
logic [384-1:0] n_s_2_00;
logic [197-1:0] n_s_0_18;
`SHADD_6(384, n_s_0_00,   0,  46,  95,  99, 103, 105, {384'b0, in0[0+:384]}, {384'b0, in0[0+:338]}, {384'b0, in0[0+:289]}, {384'b0, in0[0+:285]}, {384'b0, in0[0+:281]}, {384'b0, in0[0+:279]});
`SHADD_6(267, n_s_0_06,   0,   9,  21,  23,  28,  35, {267'b0, in0[0+:267]}, {267'b0, in0[0+:258]}, {267'b0, in0[0+:246]}, {267'b0, in0[0+:244]}, {267'b0, in0[0+:239]}, {267'b0, in0[0+:232]});
`SHADD_6(229, n_s_0_12,   0,   4,  13,  23,  25,  30, {229'b0, in0[0+:229]}, {229'b0, in0[0+:225]}, {229'b0, in0[0+:216]}, {229'b0, in0[0+:206]}, {229'b0, in0[0+:204]}, {229'b0, in0[0+:199]});
`SHADD_6(197, n_s_0_18,   0,   5,  16,  20,  22,  25, {197'b0, in0[0+:197]}, {197'b0, in0[0+:192]}, {197'b0, in0[0+:181]}, {197'b0, in0[0+:177]}, {197'b0, in0[0+:175]}, {197'b0, in0[0+:172]});
`SHADD_6(166, n_s_0_24,   0,   4,   6,  13,  16,  19, {166'b0, in0[0+:166]}, {166'b0, in0[0+:162]}, {166'b0, in0[0+:160]}, {166'b0, in0[0+:153]}, {166'b0, in0[0+:150]}, {166'b0, in0[0+:147]});
`SHADD_6(136, n_s_0_30,   0,   2,   5,  10,  12,  18, {136'b0, in0[0+:136]}, {136'b0, in0[0+:134]}, {136'b0, in0[0+:131]}, {136'b0, in0[0+:126]}, {136'b0, in0[0+:124]}, {136'b0, in0[0+:118]});
`SHADD_6(107, n_s_0_36,   0,  10,  30,  35,  45,  52, {107'b0, in0[0+:107]}, {107'b0, in0[0+: 97]}, {107'b0, in0[0+: 77]}, {107'b0, in0[0+: 72]}, {107'b0, in0[0+: 62]}, {107'b0, in0[0+: 55]});
`SHADD_6( 52, n_s_0_42,   0,  10,  12,  16,  25,  43, {52'b0, in0[0+: 52]}, {52'b0, in0[0+: 42]}, {52'b0, in0[0+: 40]}, {52'b0, in0[0+: 36]}, {52'b0, in0[0+: 27]}, {52'b0, in0[0+:  9]});
`SHADD_6(  2, n_s_0_48,   0,   0,   0,   0,   0,   0, {2'b0, in0[0+:  2]}, {2'b0, '0}, {2'b0, '0}, {2'b0, '0}, {2'b0, '0}, {2'b0, '0});
`SHADD_6(384, n_s_1_00,   0, 117, 155, 187, 218, 248, {384'b0, n_s_0_00}, {384'b0, n_s_0_06}, {384'b0, n_s_0_12}, {384'b0, n_s_0_18}, {384'b0, n_s_0_24}, {384'b0, n_s_0_30});
`SHADD_6(107, n_s_1_06,   0,  55, 105,   0,   0,   0, {107'b0, n_s_0_36}, {107'b0, n_s_0_42}, {107'b0, n_s_0_48}, {107'b0, '0}, {107'b0, '0}, {107'b0, '0});
`SHADD_6(384, n_s_2_00,   0, 277,   0,   0,   0,   0, {384'b0, n_s_1_00}, {384'b0, n_s_1_06}, {384'b0, '0}, {384'b0, '0}, {384'b0, '0}, {384'b0, '0});
assign out_n = n_s_2_00 << 0;
assign n_m_o = n_m_o_p[6-1];
always@(posedge clk) n_m_o_p[0] <= m_i;
always@(posedge clk) n_m_o_p[1] <= n_m_o_p[1-1];
always@(posedge clk) n_m_o_p[2] <= n_m_o_p[2-1];
always@(posedge clk) n_m_o_p[3] <= n_m_o_p[3-1];
always@(posedge clk) n_m_o_p[4] <= n_m_o_p[4-1];
always@(posedge clk) n_m_o_p[5] <= n_m_o_p[5-1];
always@(posedge clk) out0 <= out_p - out_n;
always@(posedge clk) m_o <= p_m_o;
endmodule

